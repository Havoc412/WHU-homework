`include "Define.v"

module test (
        input clk,

    );

endmodule