`include "Define.v"

module EXT( 
    input clk,

    input [4: 0]    iimm_shamt,
    input [11:0]	iimm, //instr[31:20], 12 bits
    input [11:0]	simm, //instr[31:25, 11:7], 12 bits
    input [11:0]	bimm, //instrD[31],instrD[7], instrD[30:25], instrD[11:8], 12 bits
    input [19:0]	uimm,
    input [19:0]	jimm_jal,

    input [6: 0]	extCtrl,

    output reg [31:0] immout
    );

    always @ (*) begin
        case (extCtrl)
            `EXT_CTRL_SHAMT:    immout <= { 27'b0, iimm_shamt[4: 0]};
            `EXT_CTRL_ITYPE:    immout <= { { (`XLEN-12){ iimm[11]}}, iimm[11: 0]}; // info 两种写法。
            `EXT_CTRL_STYPE:	immout <= { {20{ simm[11]}}, simm[11: 0]};
            // info U: 大立即数
            `EXT_CTRL_UTYPE:	immout <= { uimm[19: 0], 12'b0}; 
            // info B/J: 跳转类，左移一位。
            `EXT_CTRL_BTYPE:    immout <= { {19{ bimm[11]}}, bimm[11: 0], 1'b0};
            `EXT_CTRL_JAL:	    immout <= { {11{ jimm_jal[19]}}, jimm_jal[19: 0], 1'b0};

            default:  immout <= 32'b0;
        endcase
    end

endmodule