module My_Journey_Begins; 
  initial begin
    $display(" Hello World!" ) ;
  end
endmodule
