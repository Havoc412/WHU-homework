package PipeReg; // info 暂时不打算使用了
    
    // tag IF/ ID
    typedef struct packed {
        logic [8: 0] Cur_pc;
        logic [31: 0] Cur_Instr;
    } IF_ID_reg;

    // tag ID / EX
    typedef struct packed {
        logic ALU2ndOperandSrc; // question
        logic wrRegDataSrc; // question
        logic regWrite;
        logic memRead;
        logic memWrite;

        logic [1: 0] aluCtrl;
        logic branch;
        logic jalSel;   // question
        logic jaleSel;

        logic [1: 0] RWSel; // question

        logic [8: 0] Cur_pc;
        logic [31: 0] Cur_Instr;

        logic [31: 0] RD1;
        logic [31: 0] RD2;
        logic [4: 0] RS1; // question
        logic [4: 0] RS2;
        logic [4: 0] rd; // Immediate value generated by Imm_gen

        logic [31: 0] immGen;
        logic [2: 0] func3;
        logic [6: 0] func7;

    } ID_EX_reg;

    // tag EX / MEM
    typedef struct packed {
        logic regWrite;
        logic wrRegDataSrc;
        logic memRead;
        logic memWrite;
        logic [1: 0] RWSel; // question
        
        logic [31: 0] pc_imm;
        logic [31: 0] pc_four; // question

        logic [31: 0] immGen;
        logic [31: 0] aluRes;
        logic [31: 0] memWeData;

        logic [4: 0] rd;

        logic [2: 0] func3;
        logic [6: 0] func7;

        logic [31: 0] Cur_Instr;

    } EX_MEN_reg;

    // tag MEM / WB
    typedef struct packed {
        logic regWrite;
        logic wrRegDataSrc;
        logic [1: 0] RWSel;
        logic [31: 0] pc_imm;
        logic [31: 0] pc_four;
        logic [31: 0] immGen;
        logic [31: 0] aluRes;
        logic [31: 0] memReadData;

        logic [4: 0] rd;
        logic [31: 0] Cur_Instr;
    } MEM_WB_reg;

endpackage;