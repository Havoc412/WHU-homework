module Wave (
    input a,
    input b,
    input c
);

endmodule